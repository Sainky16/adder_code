module adder(input a,b, output sum);
    assign sum = a+b;
endmodule
